module HelloWorld;

  initial begin
    $display("Hello, World!");
    $finish; // Terminate simulation
  end

endmodule
